    Mac OS X            	   2   �      �                                      ATTR       �   �   >                  �   >  com.apple.quarantine q/0087;63ee8d57;WhatsApp;5BAD09DB-9D8E-4B9E-8AE4-1C413F64C443 